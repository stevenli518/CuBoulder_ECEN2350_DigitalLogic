`ifdef h2z
   
    divide_by = 5_000_000;
    
    
`else

    divide_by = 2_000_000;

    
`endif